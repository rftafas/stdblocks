library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;
  use IEEE.math_real.all;

package fifo_lib is

  type mem_t is ("block", "ultra", "registers", "distributed");
  attribute ram_style : string;


end package;

package body fifo_lib is



end package body;
