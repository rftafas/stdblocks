library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;
  use IEEE.math_real.all;
library expert;
  use expert.std_logic_expert.all;
library stdblocks;
    use stdblocks.ram_lib.all;

package fifo_lib is

  type fifo_status is record
    overflow  : std_logic;
    full      : std_logic;
    gofull    : std_logic;
    steady    : std_logic;
    goempty   : std_logic;
    empty     : std_logic;
    underflow : std_logic;
  end record fifo_status;

  type fifo_t is (blockram, ultra, registers, distributed);
  function fifo_type_dec ( ram_type : fifo_t ) return mem_t;

  type fifo_state_t is (underflow_st, empty_st, goempty_st, steady_st, gofull_st, full_st, overflow_st);
  function sync_state (
    ien : std_logic; oen : std_logic; iaddr : std_logic_vector; oaddr : std_logic_vector; current_state : fifo_state_t
  ) return fifo_state_t;

  function async_state (
    ien : std_logic; oen : std_logic; iaddr : std_logic_vector; oaddr : std_logic_vector; current_state : fifo_state_t
  ) return fifo_state_t;

  component stdfifo2ck
    generic (
      ram_type  : fifo_t := blockram;
      fifo_size : integer := 8;
      port_size : integer := 8
    );
    port (
      clka_i          : in  std_logic;
      rsta_i          : in  std_logic;
      clkb_i          : in  std_logic;
      rstb_i          : in  std_logic;
      dataa_i         : in  std_logic_vector(port_size-1 downto 0);
      datab_o         : out std_logic_vector(port_size-1 downto 0);
      ena_i           : in  std_logic;
      enb_i           : in  std_logic;
      fifo_status_a_o : out fifo_status;
      fifo_status_b_o : out fifo_status
    );
  end component stdfifo2ck;

  component stdfifo1ck
    generic (
      ram_type  : fifo_t := blockram;
      port_size : integer := 8;
      fifo_size : integer := 8
    );
    port (
      clk_i         : in  std_logic;
      rst_i         : in  std_logic;
      dataa_i       : in  std_logic_vector(port_size-1 downto 0);
      datab_o       : out std_logic_vector(port_size-1 downto 0);
      ena_i         : in  std_logic;
      enb_i         : in  std_logic;
      fifo_status_o : out fifo_status
    );
  end component stdfifo1ck;

  component srfifo1ck
    generic (
      fifo_size : integer := 8;
      port_size : integer := 8
    );
    port (
      clk_i         : in  std_logic;
      rst_i         : in  std_logic;
      dataa_i       : in  std_logic_vector(port_size-1 downto 0);
      datab_o       : out std_logic_vector(port_size-1 downto 0);
      ena_i         : in  std_logic;
      enb_i         : in  std_logic;
      fifo_status_o : out fifo_status
    );
  end component srfifo1ck;

  --axi parameters
  type fifo_data_rec is record
    tdest  : std_logic_vector;
    tdata  : std_logic_vector;
    tuser  : std_logic_vector;
    tlast  : std_logic;
  end record;

  type fifo_config_rec is record
    ram_type     :  fifo_t;
    fifo_size    : integer;
    tdata_size   : integer;
    tdest_size   : integer;
    tuser_size   : integer;
    packet_mode  : boolean;
    tuser_enable : boolean;
    tdest_enable : boolean;
    tlast_enable : boolean;
    cut_through  : boolean;
    sync_mode    : boolean;
  end record;

end package;

package body fifo_lib is

  function fifo_type_dec ( ram_type : fifo_t ) return mem_t is
      --variable tmp : string;
  begin
      case ram_type is
          when blockram =>
              return blockram;
          when ultra =>
              return ultra;
          when registers =>
              return registers;
          when distributed =>
              return distributed;
          when others =>
              return registers;
              report "Unknown fifo type. Using Flip-flops." severity warning;
      end case;
      --return tmp;
  end function fifo_type_dec;


  function sync_state (
    ien : std_logic; oen : std_logic; iaddr : std_logic_vector; oaddr : std_logic_vector; current_state : fifo_state_t
  ) return fifo_state_t is
    variable tmp         : fifo_state_t := steady_st;
    variable delta       : unsigned(iaddr'range) := (others=>'0');
    variable up          : std_logic             := '0';
    variable dn          : std_logic             := '0';
    variable fifo_length : integer               := 2**iaddr'length;
  begin
    tmp   := current_state;
    delta := unsigned(iaddr - oaddr);

    up := ien and not oen;
    dn := oen and not ien;

		case current_state is
      when empty_st =>
        if dn = '1' then
          tmp := underflow_st;
        elsif up = '1' then
          tmp:= goempty_st;
        end if;

      when goempty_st =>
        if delta = 1 and dn  = '1' then
          tmp :=  empty_st;
        elsif delta = fifo_length/4 then
          tmp:= steady_st;
        end if;

      when steady_st =>
        if    delta =  fifo_length/4-1 then
          tmp := goempty_st;
        elsif delta = 3*fifo_length/4 then
          tmp:= gofull_st;
        end if;

      when gofull_st =>
        if delta = fifo_length-1 and up = '1' then
          tmp:= full_st;
        elsif delta = 3*fifo_length/4-1 then
          tmp :=  steady_st;
        end if;

      when full_st =>
        if up = '1' then
          tmp :=  overflow_st;
        elsif dn = '1' then
          tmp := gofull_st;
        end if;

      when overflow_st =>
        if delta = 3*fifo_length/4-1 then
          tmp :=  steady_st;
        end if;

      when underflow_st =>
        if delta = fifo_length/4 then
          tmp:= steady_st;
        end if;

      when others =>
        tmp := steady_st;

    end case;
    return tmp;
	end sync_state;

  function async_state (
    ien : std_logic; oen : std_logic; iaddr : std_logic_vector; oaddr : std_logic_vector; current_state : fifo_state_t
  ) return fifo_state_t is
    variable tmp         : fifo_state_t := steady_st;
    variable delta       : unsigned(iaddr'range) := (others=>'0');
    variable fifo_length : integer               := 2**iaddr'length;
  begin
    tmp   := current_state;
    delta := unsigned(iaddr - oaddr);

		case current_state is

      when underflow_st =>
        if delta = fifo_length/4 then
          tmp:= steady_st;
        end if;

      when empty_st =>
        if oen = '1' then
          tmp := underflow_st;
        elsif delta = 1 then
          tmp:= goempty_st;
        end if;

      when goempty_st =>
        if delta = 1 and oen = '1' then
          tmp :=  empty_st;
        elsif delta = 0 then
          tmp :=  empty_st;
        elsif delta = fifo_length/4 then
          tmp:= steady_st;
        end if;

      when steady_st =>
        if delta = fifo_length/4-1 then
          tmp := goempty_st;
        elsif delta = 3*fifo_length/4 then
          tmp:= gofull_st;
        end if;

      when gofull_st =>
        if delta = fifo_length-1 and ien = '1' then
          tmp:= full_st;
        elsif delta = 0 then --estourou o contador.
            tmp:= full_st;
        elsif delta = 3*fifo_length/4-1 then
          tmp :=  steady_st;
        end if;

      when full_st =>
        if ien = '1' then
          tmp :=  overflow_st;
        elsif delta = fifo_length - 1 then
          tmp := gofull_st;
        end if;

      when overflow_st =>
        if delta = 3*fifo_length/4-1 then
          tmp :=  steady_st;
        end if;

      when others =>
        tmp := steady_st;

    end case;
    return tmp;
	end async_state;

---------------------------------------------------------------------------------------------------------
  function header_size_f (
    param   : fifo_config_rec
  )
  return integer is
      variable tmp : integer;
  begin
    tmp := 0;
    if not param.packet_mode then
      if param.tlast_enable then
        tmp := 1;
      end if;
      if param.tuser_enable then
        tmp := param.tuser_size + tmp;
      end if;
      if param.tdest_enable then
        tmp := tmp + param.tdest_size;
      end if;
    end if;
    return tmp;
  end header_size_f;

  function fifo_size_f (
    param   : fifo_config_rec
  )
  return integer is
      variable tmp : integer;
  begin
    tmp := param.tdata_size;
    if not param.packet_mode then
      tmp := tmp + header_size_f(param);
    end if;
    return tmp;
  end fifo_size_f;

  procedure data_bus_in (
    signal data      : in fifo_data_rec;
    param            : in fifo_config_rec;
    signal fifo_data : out std_logic_vector;
    signal head_data : out std_logic_vector
  ) is
    variable head_data_v : std_logic_vector(header_size_f(param) downto 0);
  begin
  --
    if param.tuser_enable then
      head_data_v := head_data_v sll param.tuser_size;
      head_data_v(data.tuser'range) := data.tuser;
    end if;
    if param.tdest_enable then
      head_data_v := head_data_v sll param.tdest_size;
      head_data_v(data.tdest'range) := data.tdest;
    end if;

    if param.packet_mode or param.tlast_enable then
      if param.packet_mode then
        head_data <= head_data_v;
        fifo_data <= data.tlast & data.tdata;
      else
        head_data <= (others=>'0');
        fifo_data <= data.tlast & head_data_v & data.tdata;
      end if; 
    else
      if param.packet_mode then
        head_data <= head_data_v;
        fifo_data <= data.tdata;
      else
        head_data <= (others=>'0');
        fifo_data <= head_data_v & data.tdata;
      end if;
    end if;
  end data_bus_in;

  procedure data_bus_out (
    signal data      : out fifo_data_rec;
    param            : in  fifo_config_rec;
    signal fifo_data : in  std_logic_vector;
    signal head_data : in  std_logic_vector
  ) is
    variable head_data_v : std_logic_vector(header_size_f(param)-1 downto 0);
  begin
    data.tdata  <= (others=>'0');
    data.tdest  <= (others=>'0');
    data.tuser  <= (others=>'0');
    data.tlast  <= '0';
    head_data_v := (others=>'0');

    if param.packet_mode then
      data.tdata  <= fifo_data;
      head_data_v := head_data;
    else
      data.tdata  <= fifo_data(param.tdata_size-1 downto 0);
      head_data_v := fifo_data(fifo_data'high downto param.tdata_size);
    end if;

    if param.tdest_enable then
      data.tdest  <= head_data_v(data.tdest'range);
      head_data_v := head_data_v srl param.tdest_size;
    end if;

    if param.tuser_enable then
      data.tuser  <= head_data_v(data.tuser'range);
      head_data_v := head_data_v srl param.tuser_size;
    end if;

    if param.packet_mode or param.tlast_enable then
      data.tlast <= head_data_v(0);
    end if;

  end data_bus_out;


end package body;
